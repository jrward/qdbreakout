module blocks_pos_rom(	input clk,
						input [3:0] addr,
						output reg [18:0] q	);
						
	always @ (posedge clk)
	begin
	
	/*
	100	190	280	370	460	550	145	235
325	415	505	190	280	370	460	0
320	320	320	320	320	320	330	330
330	330	330	340	340	340	340	0 */
		case (addr)
			5'h0: q <= {10'd100,9'd320};
			5'h1: q <= {10'd190,9'd320};
			5'h2: q <= {10'd280,9'd320};
			5'h3: q <= {10'd370,9'd320};
			5'h4: q <= {10'd460,9'd320};
			5'h5: q <= {10'd550,9'd320};
			5'h6: q <= {10'd145,9'd330};
			5'h7: q <= {10'd235,9'd330};
			5'h8: q <= {10'd325,9'd330};
			5'h9: q <= {10'd415,9'd330};
			5'hA: q <= {10'd505,9'd330};
			5'hB: q <= {10'd190,9'd340};
			5'hC: q <= {10'd280,9'd340};
			5'hD: q <= {10'd370,9'd340};
			5'hE: q <= {10'd460,9'd340};
			5'hF: q <= {10'd0,9'd0};
		endcase
	end
						

endmodule

